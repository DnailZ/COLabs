
module MemSim();



dist_mem_gen_0 dict(
    
)

endmodule