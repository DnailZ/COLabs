
module RAMSim;
reg rst = 0;
BM_sim b();
DM_sim d();
endmodule
